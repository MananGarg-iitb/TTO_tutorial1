/*
 * Copyright (c) 2024 Your Name
 * SPDX-License-Identifier: Apache-2.0
 */

`default_nettype none

module tt_um_example (
    input  wire [7:0] ui_in,    // Dedicated inputs
    output wire [7:0] uo_out,   // Dedicated outputs
    input  wire [7:0] uio_in,   // IOs: Input path
    output wire [7:0] uio_out,  // IOs: Output path
    output wire [7:0] uio_oe,   // IOs: Enable path (active high: 0=input, 1=output)
    input  wire       ena,      // always 1 when the design is powered, so you can ignore it
    input  wire       clk,      // clock
    input  wire       rst_n     // reset_n - low to reset
);
    
  // All output pins must be assigned. If not used, assign to 0.
  assign uio_out = 0;
  assign uio_oe  = 0;
    assign uo_out[5:0] = 0;

  // List all unused inputs to prevent warnings
    wire _unused = &{ena, uio_in, ui_in[4:0], clk, rst_n, 1'b0};


    Full_Adder uut (.A(ui_in[7]), .B(ui_in[6]), .Cin(ui_in[5]), .S(uo_out[7]), .Cout(uo_out[6]));
endmodule

module Full_Adder(
	input A,
	input B,
	input Cin,
	output S,
	output Cout
);

assign S = (A^B)^Cin;
assign Cout = (A&B)|(B&Cin)|(Cin&A);

endmodule
